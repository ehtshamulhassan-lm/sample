//This is a random file
module rand(clk, reset);
  input clk;
  input reset;
endmodule
